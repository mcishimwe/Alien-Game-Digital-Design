CONFIGURATION disp_rst_fsm_config OF disp_rst IS
   FOR fsm
   END FOR;
END disp_rst_fsm_config;