--* ><(((('> * Puli puli * ><(((('> // Ƹ̵̡Ӝ̵̨̄Ʒ * swish swish* Ƹ̵̡Ӝ̵̨̄Ʒ Ƹ̵̡Ӝ̵̨̄Ʒ // (っ◕‿◕)╭∩╮^H^H^Hっ
LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ENTITY disp_serial_tx IS PORT(bit_in:IN std_logic;clk:IN std_logic;rst_n:IN std_logic;run:IN std_logic;ready_out:OUT std_logic;s_clk:OUT std_logic;s_sda:OUT std_logic);END disp_serial_tx ;LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ARCHITECTURE fsm OF disp_serial_tx IS SIGNAL z8c3109cee:std_logic;TYPE STATE_TYPE IS(z300f5740b,zb829a35c7,z670bdf3fb);SIGNAL zdf0be1ce6:STATE_TYPE;SIGNAL ze8e79043b:STATE_TYPE;SIGNAL zddc9dc0bc:std_logic_vector(2 DOWNTO 0);SIGNAL z28618b6b9:std_logic_vector(2 DOWNTO 0);SIGNAL za21ed1d6a:std_logic;SIGNAL z0fef2b031:std_logic;SIGNAL z3a8d7a42c:std_logic;BEGIN z9149816e0:PROCESS(clk,rst_n)BEGIN IF(rst_n='0')THEN zdf0be1ce6<=z300f5740b;zddc9dc0bc<=(OTHERS=>'0');z8c3109cee<='0';ELSIF(clk'EVENT AND clk='1')THEN zdf0be1ce6<=ze8e79043b;zddc9dc0bc<=z28618b6b9;CASE zdf0be1ce6 IS WHEN z300f5740b=>z8c3109cee<=bit_in;WHEN OTHERS=>NULL;END CASE;END IF;END PROCESS z9149816e0;z145fbcc0d:PROCESS(za21ed1d6a,zdf0be1ce6,run)BEGIN z0fef2b031<='0';z3a8d7a42c<='0';CASE zdf0be1ce6 IS WHEN z300f5740b=>IF(run='1')THEN ze8e79043b<=zb829a35c7;z0fef2b031<='1';ELSE ze8e79043b<=z300f5740b;END IF;WHEN zb829a35c7=>IF(za21ed1d6a='1')THEN ze8e79043b<=z670bdf3fb;z3a8d7a42c<='1';ELSE ze8e79043b<=zb829a35c7;END IF;WHEN z670bdf3fb=>IF(za21ed1d6a='1')THEN ze8e79043b<=z300f5740b;ELSE ze8e79043b<=z670bdf3fb;END IF;WHEN OTHERS=>ze8e79043b<=z300f5740b;END CASE;END PROCESS z145fbcc0d;z822bdb2c3:PROCESS(zdf0be1ce6,z8c3109cee)BEGIN ready_out<='0';s_clk<='0';s_sda<='0';CASE zdf0be1ce6 IS WHEN z300f5740b=>ready_out<='1';WHEN zb829a35c7=>s_sda<=z8c3109cee;WHEN z670bdf3fb=>s_clk<='1';s_sda<=z8c3109cee;WHEN OTHERS=>NULL;END CASE;END PROCESS z822bdb2c3;zc4c7d2805:PROCESS(zddc9dc0bc,z0fef2b031,z3a8d7a42c)VARIABLE z35e1a2c8c:std_logic;BEGIN IF(unsigned(zddc9dc0bc)=0)THEN z35e1a2c8c:='1';ELSE z35e1a2c8c:='0';END IF;IF(z0fef2b031='1')THEN z28618b6b9<="010";ELSIF(z3a8d7a42c='1')THEN z28618b6b9<="011";ELSE IF(z35e1a2c8c='1')THEN z28618b6b9<=(OTHERS=>'0');ELSE z28618b6b9<=unsigned(zddc9dc0bc)-'1';END IF;END IF;za21ed1d6a<=z35e1a2c8c;END PROCESS zc4c7d2805;END fsm;