CONFIGURATION disp_gamma_fsm_config OF disp_gamma IS
   FOR fsm
   END FOR;
END disp_gamma_fsm_config;