CONFIGURATION reg_bank_1px_struct_config OF reg_bank_1px IS
   FOR struct
   END FOR;
END reg_bank_1px_struct_config;