CONFIGURATION mem_ctl_block_fsm_config OF mem_ctl_block IS
   FOR fsm
   END FOR;
END mem_ctl_block_fsm_config;