CONFIGURATION disp_serial_tx_fsm_config OF disp_serial_tx IS
   FOR fsm
   END FOR;
END disp_serial_tx_fsm_config;