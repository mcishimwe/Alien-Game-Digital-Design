CONFIGURATION disp_serial_led_cannon_fsm_config OF disp_serial_led_cannon IS
   FOR fsm
   END FOR;
END disp_serial_led_cannon_fsm_config;