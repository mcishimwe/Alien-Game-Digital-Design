--
-- VHDL Entity pre_made.HELLO_ALIEN.arch_name
--
-- Created:
--          by - rpmais.UNKNOWN (HTC219-304-SPC)
--          at - 13:14:04 12.10.2024
--
-- using Mentor Graphics HDL Designer(TM) 2019.3 (Build 4)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY HELLO_ALIEN IS
   PORT( 
      btn     : IN     std_logic_vector (3 DOWNTO 0);
      clk     : IN     std_logic;
      rst_n   : IN     std_logic;
      channel : OUT    std_logic_vector (7 DOWNTO 0);
      lat     : OUT    std_logic;
      s_clk   : OUT    std_logic;
      s_rst   : OUT    std_logic;
      s_sda   : OUT    std_logic;
      sb      : OUT    std_logic
   );

-- Declarations

END HELLO_ALIEN ;


--
-- VHDL Architecture pre_made.HELLO_ALIEN.struct
--
-- Created:
--          by - rpmais.UNKNOWN (HTC219-320-SPC)
--          at - 19:32:56  4.12.2024
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2019.3 (Build 4)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

LIBRARY alien_game_lib;
LIBRARY pre_made;

ARCHITECTURE struct OF HELLO_ALIEN IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL alien_col : std_logic_vector(23 DOWNTO 0);
   SIGNAL enable    : std_logic;
   SIGNAL q         : std_logic;
   SIGNAL write     : std_logic;
   SIGNAL x_coord   : std_logic_vector(7 DOWNTO 0);
   SIGNAL y_coord   : std_logic_vector(7 DOWNTO 0);


   -- ModuleWare signal declarations(v1.12) for instance 'convenience_ff' of 'adff'
   SIGNAL mw_convenience_ffreg_cval : std_logic;

   -- Component Declarations
   COMPONENT c3_t1_basic_alien
   PORT (
      clk       : IN     std_logic ;
      enable    : IN     std_logic ;
      hit       : IN     std_logic ;
      rst_n     : IN     std_logic ;
      alien_col : OUT    std_logic_vector (23 DOWNTO 0);
      alien_def : OUT    std_logic ;
      x_coord   : OUT    std_logic_vector (7 DOWNTO 0);
      y_coord   : OUT    std_logic_vector (7 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT display_controller
   PORT (
      clk        : IN     std_logic ;
      color_BGR  : IN     std_logic_vector (23 DOWNTO 0);
      frame_done : IN     std_logic ;
      rst_n      : IN     std_logic ;
      write      : IN     std_logic ;
      x_coord    : IN     std_logic_vector (7 DOWNTO 0);
      y_coord    : IN     std_logic_vector (7 DOWNTO 0);
      channel    : OUT    std_logic_vector (7 DOWNTO 0);
      lat        : OUT    std_logic ;
      s_clk      : OUT    std_logic ;
      s_rst      : OUT    std_logic ;
      s_sda      : OUT    std_logic ;
      sb         : OUT    std_logic ;
      w_rdy      : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT en_wr
   PORT (
      clk    : IN     std_logic;
      rst_n  : IN     std_logic;
      enable : OUT    std_logic;
      wr     : OUT    std_logic
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : c3_t1_basic_alien USE ENTITY alien_game_lib.c3_t1_basic_alien;
   FOR ALL : display_controller USE ENTITY pre_made.display_controller;
   FOR ALL : en_wr USE ENTITY pre_made.en_wr;
   -- pragma synthesis_on


BEGIN

   -- ModuleWare code(v1.12) for instance 'convenience_ff' of 'adff'
   q <= mw_convenience_ffreg_cval;
   convenience_ffseq_proc: PROCESS (clk, rst_n)
   BEGIN
      IF (rst_n = '0') THEN
         mw_convenience_ffreg_cval <= '0';
      ELSIF (clk'EVENT AND clk='1') THEN
         mw_convenience_ffreg_cval <= write;
      END IF;
   END PROCESS convenience_ffseq_proc;

   -- Instance port mappings.
   U_1 : c3_t1_basic_alien
      PORT MAP (
         clk       => clk,
         enable    => enable,
         hit       => btn(0),
         rst_n     => rst_n,
         alien_col => alien_col,
         alien_def => OPEN,
         x_coord   => x_coord,
         y_coord   => y_coord
      );
   U_0 : display_controller
      PORT MAP (
         clk        => clk,
         color_BGR  => alien_col,
         frame_done => q,
         rst_n      => rst_n,
         write      => write,
         x_coord    => x_coord,
         y_coord    => y_coord,
         channel    => channel,
         lat        => lat,
         s_clk      => s_clk,
         s_rst      => s_rst,
         s_sda      => s_sda,
         sb         => sb,
         w_rdy      => OPEN
      );
   U_2 : en_wr
      PORT MAP (
         clk    => clk,
         rst_n  => rst_n,
         enable => enable,
         wr     => write
      );

END struct;
